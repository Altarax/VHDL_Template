----------------------------------------------------------------------------------
--!
--! \file main.vhd
--!
--! \brief Main file.
--!
--! \version 1.0
--! \date XX/XX/XXXX
--!
--! \author Dangremont Jayson, dangremontjayson.pro@gmail.com
--!
----------------------------------------------------------------------------------

--! Use standard librairies
library library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

--! \brief Entity of the main file
--! \details Description

entity main is
    port (

        clk         : in std_logic;
        reset       : in std_logic;

        data_out    : out std_logic
        
    );
end entity main;