library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package my_types is

        type bus_array is array(natural range <>) of std_logic_vector;

end my_types;
