----------------------------------------------------------------------------------
--!
--! \file TOP_LEVEL_tb.vhd
--!
--! \brief Testbenchs for TOP_LEVEL.
--!
--! \version 1.0
--! \date XX/XX/XX
--!
--! \author Dangremont Jayson, dangremontjayson.pro@gmail.com
--!
----------------------------------------------------------------------------------

--! Use simulation librairies
Library IEEE;
use IEEE.std_logic_TEXTIO.all;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;